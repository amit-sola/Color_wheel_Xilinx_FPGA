`timescale 1ns / 1ps

// n4fpga.v - Top level module for the ECE 544 Getting Started project
//
// 
// Created By:	Roy Kravitz
// modified By: Amit Solapurkar
// Date:		23-January-2018
// Version:		1.0
//
// Description:
// ------------
// This module provides the top level for the Getting Started hardware.
// The module assume that a PmodOLED is plugged into the JA 
// expansion ports and that a PmodENC is plugged into the JD expansion 
// port (bottom row).  
//////////////////////////////////////////////////////////////////////
module n4fpga(
    input				clk,			// 100Mhz clock input
    input				btnC,			// center pushbutton
    input				btnU,			// UP (North) pusbhbutton
    input				btnL,			// LEFT (West) pushbutton
    input				btnD,			// DOWN (South) pushbutton  - used for system reset
    input				btnR,			// RIGHT (East) pushbutton
	input				btnCpuReset,	// CPU reset pushbutton
    input	[15:0]		sw,				// slide switches on Nexys 4
    output	[15:0] 		led,			// LEDs on Nexys 4   
    output              RGB1_Blue,      // RGB1 LED (LD16) 
    output              RGB1_Green,
    output              RGB1_Red,
    output              RGB2_Blue,      // RGB2 LED (LD17)
    output              RGB2_Green,
    output              RGB2_Red,
    output [7:0]        an,             // Seven Segment display
    output [6:0]        seg,
    output              dp,             // decimal point display on the seven segment 
    
    input				uart_rtl_rxd,	// USB UART Rx and Tx on Nexys 4
    output				uart_rtl_txd,	
    
	inout   [7:0]       JA,             // JA PmodOLED connector 
	                                    // both rows are used 
    output	[7:0] 		JB,				// JB Pmod connector 
                                        // Unused. Can be used for debuggin purposes 
    output	[7:0] 		JC,				// JC Pmod connector - debug signals
										// Can be used for debug purposes
	input	[7:0]		JD				// JD Pmod connector - PmodENC signals
);

// internal variables
// Clock and Reset 
wire				sysclk;             // 
wire				sysreset_n, sysreset;

// Rotary encoder 
wire				rotary_a, rotary_b, rotary_press, rotary_sw;

// GPIO pins 
wire	[7:0]	    gpio_in;				// embsys GPIO input port
wire	[7:0]	    gpio_out;				// embsys GPIO output port

wire	[31:0]		gpio1_in1;
wire	[31:0]		gpio1_in2;
wire	[31:0]		gpio2_in1;
wire	[31:0]		gpio2_in2;
wire    [31:0]      gpio3_in1;
wire    [31:0]      gpio3_in2;

wire    clk_out3;
wire	w_clk_out3;

// OLED pins 
wire 				pmodoledrgb_out_pin1_i, pmodoledrgb_out_pin1_io, pmodoledrgb_out_pin1_o, pmodoledrgb_out_pin1_t; 
wire 				pmodoledrgb_out_pin2_i, pmodoledrgb_out_pin2_io, pmodoledrgb_out_pin2_o, pmodoledrgb_out_pin2_t; 
wire 				pmodoledrgb_out_pin3_i, pmodoledrgb_out_pin3_io, pmodoledrgb_out_pin3_o, pmodoledrgb_out_pin3_t; 
wire 				pmodoledrgb_out_pin4_i, pmodoledrgb_out_pin4_io, pmodoledrgb_out_pin4_o, pmodoledrgb_out_pin4_t; 
wire 				pmodoledrgb_out_pin7_i, pmodoledrgb_out_pin7_io, pmodoledrgb_out_pin7_o, pmodoledrgb_out_pin7_t; 
wire 				pmodoledrgb_out_pin8_i, pmodoledrgb_out_pin8_io, pmodoledrgb_out_pin8_o, pmodoledrgb_out_pin8_t; 
wire 				pmodoledrgb_out_pin9_i, pmodoledrgb_out_pin9_io, pmodoledrgb_out_pin9_o, pmodoledrgb_out_pin9_t; 
wire 				pmodoledrgb_out_pin10_i, pmodoledrgb_out_pin10_io, pmodoledrgb_out_pin10_o, pmodoledrgb_out_pin10_t;

// RGB LED 
wire                w_RGB1_Red, w_RGB1_Blue, w_RGB1_Green;

// LED pins 
wire    [15:0]      led_int;                // Nexys4IO drives these outputs

// make the connections to the GPIO port.  Most of the bits are unused in the Getting
// Started project but GPIO's provide a convenient way to get the inputs and
// outputs from logic you create to and from the Microblaze.  For example,
// you may decide that using an axi_gpio peripheral is a good way to interface
// your hardware pulse-width detect logic with the Microblaze.  Our application
// is simple.
// Wrap the RGB led output back to the application program for software pulse-width detect
assign {w_RGB1_Red, w_RGB1_Blue, w_RGB1_Green} = {RGB1_Red, RGB1_Blue, RGB1_Green};
assign gpio_in = {5'b00000, w_RGB1_Red, w_RGB1_Blue, w_RGB1_Green};
assign w_clk_out3=clk_out3;
// Drive the leds from the signal generated by the microblaze 
assign led = led_int;                   // LEDs are driven by led

// make the connections
// system-wide signals
assign sysclk = clk;
assign sysreset_n = btnCpuReset;		// The CPU reset pushbutton is asserted low.  The other pushbuttons are asserted high
										// but the microblaze for Nexys 4 expects reset to be asserted low
assign sysreset = ~sysreset_n;			// Generate a reset signal that is asserted high for any logic blocks expecting it.

// Pmod OLED connections 
assign JA[0] = pmodoledrgb_out_pin1_io;
assign JA[1] = pmodoledrgb_out_pin2_io;
assign JA[2] = pmodoledrgb_out_pin3_io;
assign JA[3] = pmodoledrgb_out_pin4_io;
assign JA[4] = pmodoledrgb_out_pin7_io;
assign JA[5] = pmodoledrgb_out_pin8_io;
assign JA[6] = pmodoledrgb_out_pin9_io;
assign JA[7] = pmodoledrgb_out_pin10_io;

// JB Connector connections can be used for debug purposes
assign JB = 8'b0000000;

// JC Connector pins can be used for debug purposes 
assign JC = 8'h00; 

// PmodENC signals
// JD - bottom row only
// Pins are assigned such that turning the knob to the right
// causes the rotary count to increment.
assign rotary_a = JD[5];
assign rotary_b = JD[4];
assign rotary_press = JD[6];
assign rotary_sw = JD[7];

// instantiate the embedded system
embsys EMBSYS
       (// PMOD OLED pins 
        .PmodOLEDrgb_out_0_pin10_i(pmodoledrgb_out_pin10_i),
	    .PmodOLEDrgb_out_0_pin10_o(pmodoledrgb_out_pin10_o),
	    .PmodOLEDrgb_out_0_pin10_t(pmodoledrgb_out_pin10_t),
	    .PmodOLEDrgb_out_0_pin1_i(pmodoledrgb_out_pin1_i),
	    .PmodOLEDrgb_out_0_pin1_o(pmodoledrgb_out_pin1_o),
	    .PmodOLEDrgb_out_0_pin1_t(pmodoledrgb_out_pin1_t),
	    .PmodOLEDrgb_out_0_pin2_i(pmodoledrgb_out_pin2_i),
	    .PmodOLEDrgb_out_0_pin2_o(pmodoledrgb_out_pin2_o),
	    .PmodOLEDrgb_out_0_pin2_t(pmodoledrgb_out_pin2_t),
	    .PmodOLEDrgb_out_0_pin3_i(pmodoledrgb_out_pin3_i),
	    .PmodOLEDrgb_out_0_pin3_o(pmodoledrgb_out_pin3_o),
	    .PmodOLEDrgb_out_0_pin3_t(pmodoledrgb_out_pin3_t),
	    .PmodOLEDrgb_out_0_pin4_i(pmodoledrgb_out_pin4_i),
	    .PmodOLEDrgb_out_0_pin4_o(pmodoledrgb_out_pin4_o),
	    .PmodOLEDrgb_out_0_pin4_t(pmodoledrgb_out_pin4_t),
	    .PmodOLEDrgb_out_0_pin7_i(pmodoledrgb_out_pin7_i),
	    .PmodOLEDrgb_out_0_pin7_o(pmodoledrgb_out_pin7_o),
	    .PmodOLEDrgb_out_0_pin7_t(pmodoledrgb_out_pin7_t),
	    .PmodOLEDrgb_out_0_pin8_i(pmodoledrgb_out_pin8_i),
	    .PmodOLEDrgb_out_0_pin8_o(pmodoledrgb_out_pin8_o),
	    .PmodOLEDrgb_out_0_pin8_t(pmodoledrgb_out_pin8_t),
	    .PmodOLEDrgb_out_0_pin9_i(pmodoledrgb_out_pin9_i),
	    .PmodOLEDrgb_out_0_pin9_o(pmodoledrgb_out_pin9_o),
	    .PmodOLEDrgb_out_0_pin9_t(pmodoledrgb_out_pin9_t),
	    // GPIO pins 
        .gpio_0_GPIO_tri_i(gpio_in),
        .gpio_0_GPIO2_tri_o(gpio_out),
		.gpio_1_GPIO_tri_i(gpio1_in1),
        .gpio_1_GPIO2_tri_i(gpio1_in2),
        .gpio_2_GPIO_tri_i(gpio2_in1),
        .gpio_2_GPIO2_tri_i(gpio2_in2),
        .gpio_3_GPIO_tri_i(gpio3_in1),
        .gpio_3_GPIO2_tri_i(gpio3_in2),
        // Pmod Rotary Encoder
	    .pmodENC_A_0(rotary_a),
        .pmodENC_B_0(rotary_b),
        .pmodENC_btn_0(rotary_press),
        .pmodENC_sw_0(rotary_sw),
        // RGB1/2 Led's 
        .RGB1_Blue_0(RGB1_Blue),
        .RGB1_Green_0(RGB1_Green),
        .RGB1_Red_0(RGB1_Red),
        .RGB2_Blue_0(RGB2_Blue),
        .RGB2_Green_0(RGB2_Green),
        .RGB2_Red_0(RGB2_Red),
        // Seven Segment Display anode control  
        .an_0(an),
        .dp_0(dp),
        .led_0(led_int),
        .seg_0(seg),
        // Push buttons and switches  
        .btnC_0(btnC),
        .btnD_0(btnD),
        .btnL_0(btnL),
        .btnR_0(btnR),
        .btnU_0(btnU),
        .sw_0(sw),
        // reset and clock 
        .sysreset_n(sysreset_n),
        .sysclk(sysclk),
		.clk_out3_0(clk_out3),
        // UART pins 
        .uart_rtl_0_rxd(uart_rtl_rxd),
        .uart_rtl_0_txd(uart_rtl_txd));
  
  // Instantiating the PWM module
pwmhw pwmmodule1(w_clk_out3,w_RGB1_Red,w_RGB1_Green,w_RGB1_Blue,gpio1_in1,gpio1_in2,gpio2_in1,gpio2_in2,gpio3_in1,gpio3_in2);  
// Tristate buffers for the pmodOLEDrgb pins
// generated by PMOD bridge component.  Many
// of these signals are not tri-state.
IOBUF pmodoledrgb_out_pin1_iobuf
(
    .I(pmodoledrgb_out_pin1_o),
    .IO(pmodoledrgb_out_pin1_io),
    .O(pmodoledrgb_out_pin1_i),
    .T(pmodoledrgb_out_pin1_t)
);

IOBUF pmodoledrgb_out_pin2_iobuf
(
    .I(pmodoledrgb_out_pin2_o),
    .IO(pmodoledrgb_out_pin2_io),
    .O(pmodoledrgb_out_pin2_i),
    .T(pmodoledrgb_out_pin2_t)
);

IOBUF pmodoledrgb_out_pin3_iobuf
(
    .I(pmodoledrgb_out_pin3_o),
    .IO(pmodoledrgb_out_pin3_io),
    .O(pmodoledrgb_out_pin3_i),
    .T(pmodoledrgb_out_pin3_t)
);

IOBUF pmodoledrgb_out_pin4_iobuf
(
    .I(pmodoledrgb_out_pin4_o),
    .IO(pmodoledrgb_out_pin4_io),
    .O(pmodoledrgb_out_pin4_i),
    .T(pmodoledrgb_out_pin4_t)
);

IOBUF pmodoledrgb_out_pin7_iobuf
(
    .I(pmodoledrgb_out_pin7_o),
    .IO(pmodoledrgb_out_pin7_io),
    .O(pmodoledrgb_out_pin7_i),
    .T(pmodoledrgb_out_pin7_t)
);

IOBUF pmodoledrgb_out_pin8_iobuf
(
    .I(pmodoledrgb_out_pin8_o),
    .IO(pmodoledrgb_out_pin8_io),
    .O(pmodoledrgb_out_pin8_i),
    .T(pmodoledrgb_out_pin8_t)
);

IOBUF pmodoledrgb_out_pin9_iobuf
(
    .I(pmodoledrgb_out_pin9_o),
    .IO(pmodoledrgb_out_pin9_io),
    .O(pmodoledrgb_out_pin9_i),
    .T(pmodoledrgb_out_pin9_t)
);

IOBUF pmodoledrgb_out_pin10_iobuf
(
    .I(pmodoledrgb_out_pin10_o),
    .IO(pmodoledrgb_out_pin10_io),
    .O(pmodoledrgb_out_pin10_i),
    .T(pmodoledrgb_out_pin10_t)
);


endmodule

// PWM detection module in Hardware
module pwmhw(
input clk,
input red,
input green,
input blue,
output reg [31:0] cnt_red_high,
output reg [31:0] cnt_red_low,
output reg [31:0] cnt_green_high,
output reg [31:0] cnt_green_low,
output reg [31:0] cnt_blue_high,
output reg [31:0] cnt_blue_low

    );
     
     reg [31:0] hw_low_red = 32'd00000000;
     reg [31:0] hw_high_red = 32'd00000000;
     reg [31:0] hw_low_green = 32'd00000000;
     reg [31:0] hw_high_green = 32'd00000000;
     reg [31:0] hw_low_blue = 32'd00000000;
     reg [31:0] hw_high_blue = 32'd00000000;
     reg [31:0] timer_counter=32'd00000000;
     
     //temporary counts
     reg [31:0]           temp_red_high=32'd0;
     reg [31:0]            temp_red_low=32'd0;
     reg [31:0]           temp_green_high=32'd0;
     reg [31:0]           temp_green_low=32'd0;
     reg [31:0]             temp_blue_high=32'd0;
     reg [31:0]             temp_blue_low=32'd0;
     
     //high,low count signals
     reg [31:0]            red_high_cnt_sig=32'd0;
     reg [31:0]             red_low_cnt_sig=32'd0;
     reg [31:0]             green_high_cnt_sig=32'd0;
     reg [31:0]             green_low_cnt_sig=32'd0;
     reg [31:0]             blue_high_cnt_sig=32'd0;
     reg [31:0]             blue_low_cnt_sig=32'd0;
     
    
always @(posedge clk)
     begin
     
     //timer counter is used to adjust the frequency  e high low counts is sent to embsys module
     
     timer_counter=timer_counter+1;
     
         if(timer_counter > 32'd2)
         begin
     
         timer_counter=32'd2;
         cnt_red_high = hw_high_red;
         cnt_red_low = hw_low_red;
         cnt_green_high = hw_high_green;
         cnt_green_low = hw_low_green;
         cnt_blue_high = hw_high_blue;
         cnt_blue_low =hw_low_blue;
     
         end
     
      // Actual PWM detection Module
      // Detect Red
     
            if (red==1)
                begin
                  // Check high and low count signals
     
                  if(red_high_cnt_sig == 1 && red_low_cnt_sig == 1)
                  begin
                      hw_high_red= temp_red_high;
                      hw_low_red= temp_red_low;
     
                      temp_red_high = 1;
                      temp_red_low = 0;
     
                      red_high_cnt_sig = 0;
                      red_low_cnt_sig = 0;
     
                  end
     
                  // Increment high count
                  else
                  begin
                      red_high_cnt_sig = 1;
                      temp_red_high= temp_red_high + 1;
                  end
              end
     
              else
              begin
                  // Increment low count
                  if(red_high_cnt_sig == 1)
                  begin
                      red_low_cnt_sig = 1;
                      temp_red_low = temp_red_low + 1;
                  end
     
                  else
                       begin red_low_cnt_sig = 0; end
     
     
              end
     
              // Detect Green
     
              if(green==1)
                  begin
                      if(green_high_cnt_sig == 1 && green_low_cnt_sig == 1)
                      begin
                          hw_high_green= temp_green_high;
                          hw_low_green= temp_green_low;
     
                          temp_green_high = 1;
                          temp_green_low = 0;
     
                          green_high_cnt_sig = 0;
                          green_low_cnt_sig = 0;
     
                      end
     
                      // Increment high count
                      else
                      begin
                          green_high_cnt_sig = 1;
                          temp_green_high= temp_green_high + 1;
                      end
                  end
     
                  else
                  begin
                      // Increment low count
                      if(green_high_cnt_sig == 1)
                      begin
                          green_low_cnt_sig = 1;
                          temp_green_low = temp_green_low + 1;
                      end
     
                      else
                          green_low_cnt_sig = 0;
     
             end
     
              // Detect Blue
     
              if(blue==1)
                      begin
                          if(blue_high_cnt_sig == 1 && blue_low_cnt_sig == 1)
                          begin
                              hw_high_blue= temp_blue_high;
                              hw_low_blue= temp_blue_low;
     
                              temp_blue_high = 1;
                              temp_blue_low = 0;
     
                              blue_high_cnt_sig = 0;
                              blue_low_cnt_sig = 0;
     
                          end
     
                          // Increment high count
                          else
                          begin
                              blue_high_cnt_sig = 1;
                              temp_blue_high = temp_blue_high + 1;
                          end
                      end
     
                      else
                      begin
                          // Increment low count value
                          if(blue_high_cnt_sig == 1)
                          begin
                              blue_low_cnt_sig = 1;
                              temp_blue_low = temp_blue_low + 1;
                          end
     
                          else
                               begin blue_low_cnt_sig = 0; end
                               
                           end
          end
endmodule